`timescale 1ns/100ps
module fft_fc_layer(
	input clock,reset,
	input

	output 
	);

endmodule